module FSM (Clock,Reset);
//init


//Behavioral Verilog
reg [36:0]State;

always @ (posedge Clock) begin
	case (1'b1)
		State[0]:
		State[1]:
		State[2]:
		State[3]:
		State[4]:
		State[5]:
		State[6]:
		State[7]:
		State[8]:
		State[9]:
		State[10]:
		State[11]:
		State[12]:
		State[13]:
		State[14]:
		State[15]:
		State[16]:
		State[17]:
		State[18]:
		State[19]:
		State[20]:
		State[21]:
		State[22]:
		State[23]:
		State[24]:
		State[25]:
		State[26]:
		State[27]:
		State[28]:
		State[29]:
		State[30]:
		State[31]:
		State[32]:
		State[33]:
		State[34]:
		State[35]:

end
endmodule